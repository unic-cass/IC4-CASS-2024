VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO SLOPEDETECT
  CLASS BLOCK ;
  FOREIGN SLOPEDETECT ;
  ORIGIN 0.000 0.000 ;
  SIZE 1810.000 BY 980.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 1806.000 49.000 1810.000 49.600 ;
    END
  END io_in[0]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 1806.000 342.760 1810.000 343.360 ;
    END
  END io_in[1]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1806.000 244.840 1810.000 245.440 ;
    END
  END io_oeb[0]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1806.000 538.600 1810.000 539.200 ;
    END
  END io_oeb[1]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1806.000 734.440 1810.000 735.040 ;
    END
  END io_oeb[2]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1806.000 930.280 1810.000 930.880 ;
    END
  END io_oeb[3]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 1806.000 146.920 1810.000 147.520 ;
    END
  END io_out[0]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 1806.000 440.680 1810.000 441.280 ;
    END
  END io_out[1]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 1806.000 636.520 1810.000 637.120 ;
    END
  END io_out[2]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 1806.000 832.360 1810.000 832.960 ;
    END
  END io_out[3]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 968.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 968.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 968.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 968.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 968.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 968.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 968.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 968.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 968.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1403.440 10.640 1405.040 968.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1557.040 10.640 1558.640 968.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1710.640 10.640 1712.240 968.560 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 968.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 968.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 968.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 968.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 968.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 968.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 968.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 968.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1326.640 10.640 1328.240 968.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1480.240 10.640 1481.840 968.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1633.840 10.640 1635.440 968.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1787.440 10.640 1789.040 968.560 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 452.270 0.000 452.550 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 1357.090 0.000 1357.370 4.000 ;
    END
  END wb_rst_i
  OBS
      LAYER nwell ;
        RECT 5.330 964.185 1804.310 967.015 ;
        RECT 5.330 958.745 1804.310 961.575 ;
        RECT 5.330 953.305 1804.310 956.135 ;
        RECT 5.330 947.865 1804.310 950.695 ;
        RECT 5.330 942.425 1804.310 945.255 ;
        RECT 5.330 936.985 1804.310 939.815 ;
        RECT 5.330 931.545 1804.310 934.375 ;
        RECT 5.330 926.105 1804.310 928.935 ;
        RECT 5.330 920.665 1804.310 923.495 ;
        RECT 5.330 915.225 1804.310 918.055 ;
        RECT 5.330 909.785 1804.310 912.615 ;
        RECT 5.330 904.345 1804.310 907.175 ;
        RECT 5.330 898.905 1804.310 901.735 ;
        RECT 5.330 893.465 1804.310 896.295 ;
        RECT 5.330 888.025 1804.310 890.855 ;
        RECT 5.330 882.585 1804.310 885.415 ;
        RECT 5.330 877.145 1804.310 879.975 ;
        RECT 5.330 871.705 1804.310 874.535 ;
        RECT 5.330 866.265 1804.310 869.095 ;
        RECT 5.330 860.825 1804.310 863.655 ;
        RECT 5.330 855.385 1804.310 858.215 ;
        RECT 5.330 849.945 1804.310 852.775 ;
        RECT 5.330 844.505 1804.310 847.335 ;
        RECT 5.330 839.065 1804.310 841.895 ;
        RECT 5.330 833.625 1804.310 836.455 ;
        RECT 5.330 828.185 1804.310 831.015 ;
        RECT 5.330 822.745 1804.310 825.575 ;
        RECT 5.330 817.305 1804.310 820.135 ;
        RECT 5.330 811.865 1804.310 814.695 ;
        RECT 5.330 806.425 1804.310 809.255 ;
        RECT 5.330 800.985 1804.310 803.815 ;
        RECT 5.330 795.545 1804.310 798.375 ;
        RECT 5.330 790.105 1804.310 792.935 ;
        RECT 5.330 784.665 1804.310 787.495 ;
        RECT 5.330 779.225 1804.310 782.055 ;
        RECT 5.330 773.785 1804.310 776.615 ;
        RECT 5.330 768.345 1804.310 771.175 ;
        RECT 5.330 762.905 1804.310 765.735 ;
        RECT 5.330 757.465 1804.310 760.295 ;
        RECT 5.330 752.025 1804.310 754.855 ;
        RECT 5.330 746.585 1804.310 749.415 ;
        RECT 5.330 741.145 1804.310 743.975 ;
        RECT 5.330 735.705 1804.310 738.535 ;
        RECT 5.330 730.265 1804.310 733.095 ;
        RECT 5.330 724.825 1804.310 727.655 ;
        RECT 5.330 719.385 1804.310 722.215 ;
        RECT 5.330 713.945 1804.310 716.775 ;
        RECT 5.330 708.505 1804.310 711.335 ;
        RECT 5.330 703.065 1804.310 705.895 ;
        RECT 5.330 697.625 1804.310 700.455 ;
        RECT 5.330 692.185 1804.310 695.015 ;
        RECT 5.330 686.745 1804.310 689.575 ;
        RECT 5.330 681.305 1804.310 684.135 ;
        RECT 5.330 675.865 1804.310 678.695 ;
        RECT 5.330 670.425 1804.310 673.255 ;
        RECT 5.330 664.985 1804.310 667.815 ;
        RECT 5.330 659.545 1804.310 662.375 ;
        RECT 5.330 654.105 1804.310 656.935 ;
        RECT 5.330 648.665 1804.310 651.495 ;
        RECT 5.330 643.225 1804.310 646.055 ;
        RECT 5.330 637.785 1804.310 640.615 ;
        RECT 5.330 632.345 1804.310 635.175 ;
        RECT 5.330 626.905 1804.310 629.735 ;
        RECT 5.330 621.465 1804.310 624.295 ;
        RECT 5.330 616.025 1804.310 618.855 ;
        RECT 5.330 610.585 1804.310 613.415 ;
        RECT 5.330 605.145 1804.310 607.975 ;
        RECT 5.330 599.705 1804.310 602.535 ;
        RECT 5.330 594.265 1804.310 597.095 ;
        RECT 5.330 588.825 1804.310 591.655 ;
        RECT 5.330 583.385 1804.310 586.215 ;
        RECT 5.330 577.945 1804.310 580.775 ;
        RECT 5.330 572.505 1804.310 575.335 ;
        RECT 5.330 567.065 1804.310 569.895 ;
        RECT 5.330 561.625 1804.310 564.455 ;
        RECT 5.330 556.185 1804.310 559.015 ;
        RECT 5.330 550.745 1804.310 553.575 ;
        RECT 5.330 545.305 1804.310 548.135 ;
        RECT 5.330 539.865 1804.310 542.695 ;
        RECT 5.330 534.425 1804.310 537.255 ;
        RECT 5.330 528.985 1804.310 531.815 ;
        RECT 5.330 523.545 1804.310 526.375 ;
        RECT 5.330 518.105 1804.310 520.935 ;
        RECT 5.330 512.665 1804.310 515.495 ;
        RECT 5.330 507.225 1804.310 510.055 ;
        RECT 5.330 501.785 1804.310 504.615 ;
        RECT 5.330 496.345 1804.310 499.175 ;
        RECT 5.330 490.905 1804.310 493.735 ;
        RECT 5.330 485.465 1804.310 488.295 ;
        RECT 5.330 480.025 1804.310 482.855 ;
        RECT 5.330 474.585 1804.310 477.415 ;
        RECT 5.330 469.145 1804.310 471.975 ;
        RECT 5.330 463.705 1804.310 466.535 ;
        RECT 5.330 458.265 1804.310 461.095 ;
        RECT 5.330 452.825 1804.310 455.655 ;
        RECT 5.330 447.385 1804.310 450.215 ;
        RECT 5.330 441.945 1804.310 444.775 ;
        RECT 5.330 436.505 1804.310 439.335 ;
        RECT 5.330 431.065 1804.310 433.895 ;
        RECT 5.330 425.625 1804.310 428.455 ;
        RECT 5.330 420.185 1804.310 423.015 ;
        RECT 5.330 414.745 1804.310 417.575 ;
        RECT 5.330 409.305 1804.310 412.135 ;
        RECT 5.330 403.865 1804.310 406.695 ;
        RECT 5.330 398.425 1804.310 401.255 ;
        RECT 5.330 392.985 1804.310 395.815 ;
        RECT 5.330 387.545 1804.310 390.375 ;
        RECT 5.330 382.105 1804.310 384.935 ;
        RECT 5.330 376.665 1804.310 379.495 ;
        RECT 5.330 371.225 1804.310 374.055 ;
        RECT 5.330 365.785 1804.310 368.615 ;
        RECT 5.330 360.345 1804.310 363.175 ;
        RECT 5.330 354.905 1804.310 357.735 ;
        RECT 5.330 349.465 1804.310 352.295 ;
        RECT 5.330 344.025 1804.310 346.855 ;
        RECT 5.330 338.585 1804.310 341.415 ;
        RECT 5.330 333.145 1804.310 335.975 ;
        RECT 5.330 327.705 1804.310 330.535 ;
        RECT 5.330 322.265 1804.310 325.095 ;
        RECT 5.330 316.825 1804.310 319.655 ;
        RECT 5.330 311.385 1804.310 314.215 ;
        RECT 5.330 305.945 1804.310 308.775 ;
        RECT 5.330 300.505 1804.310 303.335 ;
        RECT 5.330 295.065 1804.310 297.895 ;
        RECT 5.330 289.625 1804.310 292.455 ;
        RECT 5.330 284.185 1804.310 287.015 ;
        RECT 5.330 278.745 1804.310 281.575 ;
        RECT 5.330 273.305 1804.310 276.135 ;
        RECT 5.330 267.865 1804.310 270.695 ;
        RECT 5.330 262.425 1804.310 265.255 ;
        RECT 5.330 256.985 1804.310 259.815 ;
        RECT 5.330 251.545 1804.310 254.375 ;
        RECT 5.330 246.105 1804.310 248.935 ;
        RECT 5.330 240.665 1804.310 243.495 ;
        RECT 5.330 235.225 1804.310 238.055 ;
        RECT 5.330 229.785 1804.310 232.615 ;
        RECT 5.330 224.345 1804.310 227.175 ;
        RECT 5.330 218.905 1804.310 221.735 ;
        RECT 5.330 213.465 1804.310 216.295 ;
        RECT 5.330 208.025 1804.310 210.855 ;
        RECT 5.330 202.585 1804.310 205.415 ;
        RECT 5.330 197.145 1804.310 199.975 ;
        RECT 5.330 191.705 1804.310 194.535 ;
        RECT 5.330 186.265 1804.310 189.095 ;
        RECT 5.330 180.825 1804.310 183.655 ;
        RECT 5.330 175.385 1804.310 178.215 ;
        RECT 5.330 169.945 1804.310 172.775 ;
        RECT 5.330 164.505 1804.310 167.335 ;
        RECT 5.330 159.065 1804.310 161.895 ;
        RECT 5.330 153.625 1804.310 156.455 ;
        RECT 5.330 148.185 1804.310 151.015 ;
        RECT 5.330 142.745 1804.310 145.575 ;
        RECT 5.330 137.305 1804.310 140.135 ;
        RECT 5.330 131.865 1804.310 134.695 ;
        RECT 5.330 126.425 1804.310 129.255 ;
        RECT 5.330 120.985 1804.310 123.815 ;
        RECT 5.330 115.545 1804.310 118.375 ;
        RECT 5.330 110.105 1804.310 112.935 ;
        RECT 5.330 104.665 1804.310 107.495 ;
        RECT 5.330 99.225 1804.310 102.055 ;
        RECT 5.330 93.785 1804.310 96.615 ;
        RECT 5.330 88.345 1804.310 91.175 ;
        RECT 5.330 82.905 1804.310 85.735 ;
        RECT 5.330 77.465 1804.310 80.295 ;
        RECT 5.330 72.025 1804.310 74.855 ;
        RECT 5.330 66.585 1804.310 69.415 ;
        RECT 5.330 61.145 1804.310 63.975 ;
        RECT 5.330 55.705 1804.310 58.535 ;
        RECT 5.330 50.265 1804.310 53.095 ;
        RECT 5.330 44.825 1804.310 47.655 ;
        RECT 5.330 39.385 1804.310 42.215 ;
        RECT 5.330 33.945 1804.310 36.775 ;
        RECT 5.330 28.505 1804.310 31.335 ;
        RECT 5.330 23.065 1804.310 25.895 ;
        RECT 5.330 17.625 1804.310 20.455 ;
        RECT 5.330 12.185 1804.310 15.015 ;
      LAYER li1 ;
        RECT 5.520 10.795 1804.120 968.405 ;
      LAYER met1 ;
        RECT 5.520 10.640 1804.420 968.560 ;
      LAYER met2 ;
        RECT 21.070 4.280 1804.030 968.505 ;
        RECT 21.070 4.000 451.990 4.280 ;
        RECT 452.830 4.000 1356.810 4.280 ;
        RECT 1357.650 4.000 1804.030 4.280 ;
      LAYER met3 ;
        RECT 21.050 931.280 1806.000 968.485 ;
        RECT 21.050 929.880 1805.600 931.280 ;
        RECT 21.050 833.360 1806.000 929.880 ;
        RECT 21.050 831.960 1805.600 833.360 ;
        RECT 21.050 735.440 1806.000 831.960 ;
        RECT 21.050 734.040 1805.600 735.440 ;
        RECT 21.050 637.520 1806.000 734.040 ;
        RECT 21.050 636.120 1805.600 637.520 ;
        RECT 21.050 539.600 1806.000 636.120 ;
        RECT 21.050 538.200 1805.600 539.600 ;
        RECT 21.050 441.680 1806.000 538.200 ;
        RECT 21.050 440.280 1805.600 441.680 ;
        RECT 21.050 343.760 1806.000 440.280 ;
        RECT 21.050 342.360 1805.600 343.760 ;
        RECT 21.050 245.840 1806.000 342.360 ;
        RECT 21.050 244.440 1805.600 245.840 ;
        RECT 21.050 147.920 1806.000 244.440 ;
        RECT 21.050 146.520 1805.600 147.920 ;
        RECT 21.050 50.000 1806.000 146.520 ;
        RECT 21.050 48.600 1805.600 50.000 ;
        RECT 21.050 10.715 1806.000 48.600 ;
      LAYER met4 ;
        RECT 232.135 150.455 251.040 817.185 ;
        RECT 253.440 150.455 327.840 817.185 ;
        RECT 330.240 150.455 404.640 817.185 ;
        RECT 407.040 150.455 481.440 817.185 ;
        RECT 483.840 150.455 558.240 817.185 ;
        RECT 560.640 150.455 635.040 817.185 ;
        RECT 637.440 150.455 711.840 817.185 ;
        RECT 714.240 150.455 788.640 817.185 ;
        RECT 791.040 150.455 865.440 817.185 ;
        RECT 867.840 150.455 942.240 817.185 ;
        RECT 944.640 150.455 1019.040 817.185 ;
        RECT 1021.440 150.455 1095.840 817.185 ;
        RECT 1098.240 150.455 1172.640 817.185 ;
        RECT 1175.040 150.455 1249.440 817.185 ;
        RECT 1251.840 150.455 1326.240 817.185 ;
        RECT 1328.640 150.455 1403.040 817.185 ;
        RECT 1405.440 150.455 1479.840 817.185 ;
        RECT 1482.240 150.455 1556.640 817.185 ;
        RECT 1559.040 150.455 1567.385 817.185 ;
  END
END SLOPEDETECT
END LIBRARY

